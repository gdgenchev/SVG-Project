<?xml version="1.0" standalone="no"?>
<!DOCTYPE svg PUBLIC "-//W3C//DTD SVG 1.1//EN" 
  "http://www.w3.org/Graphics/SVG/1.1/DTD/svg11.dtd">
<svg width="12cm" height="4cm" viewBox="0 0 1200 400"
     xmlns="http://www.w3.org/2000/svg" version="1.1">
  <desc>Example rect01 - rectangle with sharp corners</desc>

  <!-- Show outline of canvas using 'rect' element -->
  <rect x="1" y="1" width="1198" height="398"
		fill="none" stroke="blue" stroke-width="2" />

  <line x1="20" y1="100" x2="100" y2="20"
		stroke-width="2" stroke="red" />

  <rect x="20" y="30" width="40" height="50"
		fill="red" stroke="red" stroke-width="1" />

  <rect x="10" y="20" width="30" height="40"
		fill="red" stroke="blue" stroke-width="1" />

  <line x1="100" y1="200" x2="300" y2="400"
		stroke-width="2" stroke="red" />

  <circle cx="10" cy="20" r="30"
		fill="red" stroke="blue" stroke-width="2" />

</svg>
